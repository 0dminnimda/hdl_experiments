typedef buff_uart_rx_config;

