typedef buff_uart_tx_config;

