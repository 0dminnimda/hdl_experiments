class buff_uart_tx_config extends uvm_object;

