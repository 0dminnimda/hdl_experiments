class buff_uart_rx_config extends uvm_object;

